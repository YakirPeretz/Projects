// Synchronous FIFO tests package
// Create By: Yakir Peretz


package fifo_test_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    `include "YP_sync_fifo_base_tests.sv"
endpackage