// packet fifo
// Create By: Yakir Peretz

`resetall
`timescale 1ps/1ps
module InChannel_fsm #( // Parameters
parameter data_size          = 8,
parameter pkt_length_bits    = 5,
parameter pkt_addr_bits      = data_size-pkt_length_bits// 8-5 = 3
)








endmodule